`include "csa32.v"

module mult16(
    input [15:0] data1,
    input [15:0] data2,
    output [31:0] out
);

wire [15:0] p_prod [0:15]; //partial product

generate
    genvar i;
    for(i=0; i<16; i=i+1) begin
        assign p_prod[i] = data2[i] ? data1 : 16'b0;
    end    
endgenerate
wire \1/0 , \2/0 , \2/1 , \3/0 , \3/1 , \3/2 , \4/0 , \4/1 , \4/2 , \4/3 , 
    \5/0 , \5/1 , \5/2 , \5/3 , \5/4 , \6/0 , \6/1 , \6/2 , \6/3 , \6/4 , 
    \6/5 , \7/0 , \7/1 , \7/2 , \7/3 , \7/4 , \7/5 , \7/6 , \8/0 , \8/1 , 
    \8/2 , \8/3 , \8/4 , \8/5 , \8/6 , \8/7 , \9/0 , \9/1 , \9/2 , \9/3 , 
    \9/4 , \9/5 , \9/6 , \9/7 , \9/8 , \10/0 , \10/1 , \10/2 , \10/3 , \10/4 , 
    \10/5 , \10/6 , \10/7 , \10/8 , \10/9 , \11/0 , \11/1 , \11/2 , \11/3 , \11/4 , 
    \11/5 , \11/6 , \11/7 , \11/8 , \11/9 , \11/10 , \12/0 , \12/1 , \12/2 , \12/3 , 
    \12/4 , \12/5 , \12/6 , \12/7 , \12/8 , \12/9 , \12/10 , \12/11 , \13/0 , \13/1 , 
    \13/2 , \13/3 , \13/4 , \13/5 , \13/6 , \13/7 , \13/8 , \13/9 , \13/10 , \13/11 , 
    \13/12 , \14/0 , \14/1 , \14/2 , \14/3 , \14/4 , \14/5 , \14/6 , \14/7 , \14/8 , 
    \14/9 , \14/10 , \14/11 , \14/12 , \14/13 , \15/0 , \15/1 , \15/2 , \15/3 , \15/4 , 
    \15/5 , \15/6 , \15/7 , \15/8 , \15/9 , \15/10 , \15/11 , \15/12 , \15/13 , \15/14 , 
    \16/0 , \16/1 , \16/2 , \16/3 , \16/4 , \16/5 , \16/6 , \16/7 , \16/8 , \16/9 , 
    \16/10 , \16/11 , \16/12 , \16/13 , \16/14 , \16/15 , \17/0 , \17/1 , \17/2 , \17/3 , 
    \17/4 , \17/5 , \17/6 , \17/7 , \17/8 , \17/9 , \17/10 , \17/11 , \17/12 , \17/13 , 
    \17/14 , \18/0 , \18/1 , \18/2 , \18/3 , \18/4 , \18/5 , \18/6 , \18/7 , \18/8 , 
    \18/9 , \18/10 , \18/11 , \18/12 , \18/13 , \19/0 , \19/1 , \19/2 , \19/3 , \19/4 , 
    \19/5 , \19/6 , \19/7 , \19/8 , \19/9 , \19/10 , \19/11 , \19/12 , \20/0 , \20/1 , 
    \20/2 , \20/3 , \20/4 , \20/5 , \20/6 , \20/7 , \20/8 , \20/9 , \20/10 , \20/11 , 
    \21/0 , \21/1 , \21/2 , \21/3 , \21/4 , \21/5 , \21/6 , \21/7 , \21/8 , \21/9 , 
    \21/10 , \22/0 , \22/1 , \22/2 , \22/3 , \22/4 , \22/5 , \22/6 , \22/7 , \22/8 , 
    \22/9 , \23/0 , \23/1 , \23/2 , \23/3 , \23/4 , \23/5 , \23/6 , \23/7 , \23/8 , 
    \24/0 , \24/1 , \24/2 , \24/3 , \24/4 , \24/5 , \24/6 , \24/7 , \25/0 , \25/1 , 
    \25/2 , \25/3 , \25/4 , \25/5 , \25/6 , \26/0 , \26/1 , \26/2 , \26/3 , \26/4 , 
    \26/5 , \27/0 , \27/1 , \27/2 , \27/3 , \27/4 , \28/0 , \28/1 , \28/2 , \28/3 , 
    \29/0 , \29/1 , \29/2 , \30/0 , \30/1 , \31/0 , \s1 , \c1 , \s2 , \c2 , 
    \s3 , \c3 , \s4 , \c4 , \s5 , \c5 , \s6 , \c6 , \s7 , \c7 , 
    \s8 , \c8 , \s9 , \c9 , \s10 , \c10 , \s11 , \c11 , \s12 , \c12 , 
    \s13 , \c13 , \s14 , \c14 , \s15 , \c15 , \s16 , \c16 , \s17 , \c17 , 
    \s18 , \c18 , \s19 , \c19 , \s20 , \c20 , \s21 , \c21 , \s22 , \c22 , 
    \s23 , \c23 , \s24 , \c24 , \s25 , \c25 , \s26 , \c26 , \s27 , \c27 , 
    \s28 , \c28 , \s29 , \c29 , \s30 , \c30 , \s31 , \c31 , \s32 , \c32 , 
    \s33 , \c33 , \s34 , \c34 , \s35 , \c35 , \s36 , \c36 , \s37 , \c37 , 
    \s38 , \c38 , \s39 , \c39 , \s40 , \c40 , \s41 , \c41 , \s42 , \c42 , 
    \s43 , \c43 , \s44 , \c44 , \s45 , \c45 , \s46 , \c46 , \s47 , \c47 , 
    \s48 , \c48 , \s49 , \c49 , \s50 , \c50 , \s51 , \c51 , \s52 , \c52 , 
    \s53 , \c53 , \s54 , \c54 , \s55 , \c55 , \s56 , \c56 , \s57 , \c57 , 
    \s58 , \c58 , \s59 , \c59 , \s60 , \c60 , \s61 , \c61 , \s62 , \c62 , 
    \s63 , \c63 , \s64 , \c64 , \s65 , \c65 , \s66 , \c66 , \s67 , \c67 , 
    \s68 , \c68 , \s69 , \c69 , \s70 , \c70 , \s71 , \c71 , \s72 , \c72 , 
    \s73 , \c73 , \s74 , \c74 , \s75 , \c75 , \s76 , \c76 , \s77 , \c77 , 
    \s78 , \c78 , \s79 , \c79 , \s80 , \c80 , \s81 , \c81 , \s82 , \c82 , 
    \s83 , \c83 , \s84 , \c84 , \s85 , \c85 , \s86 , \c86 , \s87 , \c87 , 
    \s88 , \c88 , \s89 , \c89 , \s90 , \c90 , \s91 , \c91 , \s92 , \c92 , 
    \s93 , \c93 , \s94 , \c94 , \s95 , \c95 , \s96 , \c96 , \s97 , \c97 , 
    \s98 , \c98 , \s99 , \c99 , \s100 , \c100 , \s101 , \c101 , \s102 , \c102 , 
    \s103 , \c103 , \s104 , \c104 , \s105 , \c105 , \s106 , \c106 , \s107 , \c107 , 
    \s108 , \c108 , \s109 , \c109 , \s110 , \c110 , \s111 , \c111 , \s112 , \c112 , 
    \s113 , \c113 , \s114 , \c114 , \s115 , \c115 , \s116 , \c116 , \s117 , \c117 , 
    \s118 , \c118 , \s119 , \c119 , \s120 , \c120 , \s121 , \c121 , \s122 , \c122 , 
    \s123 , \c123 , \s124 , \c124 , \s125 , \c125 , \s126 , \c126 , \s127 , \c127 , 
    \s128 , \c128 , \s129 , \c129 , \s130 , \c130 , \s131 , \c131 , \s132 , \c132 , 
    \s133 , \c133 , \s134 , \c134 , \s135 , \c135 , \s136 , \c136 , \s137 , \c137 , 
    \s138 , \c138 , \s139 , \c139 , \s140 , \c140 , \s141 , \c141 , \s142 , \c142 , 
    \s143 , \c143 , \s144 , \c144 , \s145 , \c145 , \s146 , \c146 , \s147 , \c147 , 
    \s148 , \c148 , \s149 , \c149 , \s150 , \c150 , \s151 , \c151 , \s152 , \c152 , 
    \s153 , \c153 , \s154 , \c154 , \s155 , \c155 , \s156 , \c156 , \s157 , \c157 , 
    \s158 , \c158 , \s159 , \c159 , \s160 , \c160 , \s161 , \c161 , \s162 , \c162 , 
    \s163 , \c163 , \s164 , \c164 , \s165 , \c165 , \s166 , \c166 , \s167 , \c167 , 
    \s168 , \c168 , \s169 , \c169 , \sf1 , \cf1 , \s170 , \c170 , \s171 , \c171 , 
    \s172 , \c172 , \s173 , \c173 , \s174 , \c174 , \s175 , \c175 , \s176 , \c176 , 
    \s177 , \c177 , \s178 , \c178 , \s179 , \c179 , \s180 , \c180 , \s181 , \c181 , 
    \s182 , \c182 , \s183 , \c183 , \s184 , \c184 , \s185 , \c185 , \s186 , \c186 , 
    \s187 , \c187 , \s188 , \c188 , \s189 , \c189 , \s190 , \c190 , \s191 , \c191 , 
    \s192 , \c192 , \s193 , \c193 , \s194 , \c194 , \s195 , \c195 , \s196 , \c196 , 
    \s197 , \c197 , \s198 , \c198 , \s199 , \c199 , \s200 , \c200 , \sf2 , \cf2 , 
    \sf3 , \cf3 , \sf4 , \cf4 , \sf5 , \cf5 , \sf6 , \cf6 , \sf7 , \cf7 , 
    \sf8 , \cf8 , \sf9 , \cf9 , \s201 , \c201 , \sf10 , \cf10 ;
wire [31:0] in1, in2;
wire ov;





assign \1/0 = p_prod[15][15] ;
assign \2/0 = p_prod[14][15] ;
assign \2/1 = p_prod[15][14] ;
assign \3/0 = p_prod[13][15] ;
assign \3/1 = p_prod[14][14] ;
assign \3/2 = p_prod[15][13] ;
assign \4/0 = p_prod[12][15] ;
assign \4/1 = p_prod[13][14] ;
assign \4/2 = p_prod[14][13] ;
assign \4/3 = p_prod[15][12] ;
assign \5/0 = p_prod[11][15] ;
assign \5/1 = p_prod[12][14] ;
assign \5/2 = p_prod[13][13] ;
assign \5/3 = p_prod[14][12] ;
assign \5/4 = p_prod[15][11] ;
assign \6/0 = p_prod[10][15] ;
assign \6/1 = p_prod[11][14] ;
assign \6/2 = p_prod[12][13] ;
assign \6/3 = p_prod[13][12] ;
assign \6/4 = p_prod[14][11] ;
assign \6/5 = p_prod[15][10] ;
assign \7/0 = p_prod[9][15] ;
assign \7/1 = p_prod[10][14] ;
assign \7/2 = p_prod[11][13] ;
assign \7/3 = p_prod[12][12] ;
assign \7/4 = p_prod[13][11] ;
assign \7/5 = p_prod[14][10] ;
assign \7/6 = p_prod[15][9] ;
assign \8/0 = p_prod[8][15] ;
assign \8/1 = p_prod[9][14] ;
assign \8/2 = p_prod[10][13] ;
assign \8/3 = p_prod[11][12] ;
assign \8/4 = p_prod[12][11] ;
assign \8/5 = p_prod[13][10] ;
assign \8/6 = p_prod[14][9] ;
assign \8/7 = p_prod[15][8] ;
assign \9/0 = p_prod[7][15] ;
assign \9/1 = p_prod[8][14] ;
assign \9/2 = p_prod[9][13] ;
assign \9/3 = p_prod[10][12] ;
assign \9/4 = p_prod[11][11] ;
assign \9/5 = p_prod[12][10] ;
assign \9/6 = p_prod[13][9] ;
assign \9/7 = p_prod[14][8] ;
assign \9/8 = p_prod[15][7] ;
assign \10/0 = p_prod[6][15] ;
assign \10/1 = p_prod[7][14] ;
assign \10/2 = p_prod[8][13] ;
assign \10/3 = p_prod[9][12] ;
assign \10/4 = p_prod[10][11] ;
assign \10/5 = p_prod[11][10] ;
assign \10/6 = p_prod[12][9] ;
assign \10/7 = p_prod[13][8] ;
assign \10/8 = p_prod[14][7] ;
assign \10/9 = p_prod[15][6] ;
assign \11/0 = p_prod[5][15] ;
assign \11/1 = p_prod[6][14] ;
assign \11/2 = p_prod[7][13] ;
assign \11/3 = p_prod[8][12] ;
assign \11/4 = p_prod[9][11] ;
assign \11/5 = p_prod[10][10] ;
assign \11/6 = p_prod[11][9] ;
assign \11/7 = p_prod[12][8] ;
assign \11/8 = p_prod[13][7] ;
assign \11/9 = p_prod[14][6] ;
assign \11/10 = p_prod[15][5] ;
assign \12/0 = p_prod[4][15] ;
assign \12/1 = p_prod[5][14] ;
assign \12/2 = p_prod[6][13] ;
assign \12/3 = p_prod[7][12] ;
assign \12/4 = p_prod[8][11] ;
assign \12/5 = p_prod[9][10] ;
assign \12/6 = p_prod[10][9] ;
assign \12/7 = p_prod[11][8] ;
assign \12/8 = p_prod[12][7] ;
assign \12/9 = p_prod[13][6] ;
assign \12/10 = p_prod[14][5] ;
assign \12/11 = p_prod[15][4] ;
assign \13/0 = p_prod[3][15] ;
assign \13/1 = p_prod[4][14] ;
assign \13/2 = p_prod[5][13] ;
assign \13/3 = p_prod[6][12] ;
assign \13/4 = p_prod[7][11] ;
assign \13/5 = p_prod[8][10] ;
assign \13/6 = p_prod[9][9] ;
assign \13/7 = p_prod[10][8] ;
assign \13/8 = p_prod[11][7] ;
assign \13/9 = p_prod[12][6] ;
assign \13/10 = p_prod[13][5] ;
assign \13/11 = p_prod[14][4] ;
assign \13/12 = p_prod[15][3] ;
assign \14/0 = p_prod[2][15] ;
assign \14/1 = p_prod[3][14] ;
assign \14/2 = p_prod[4][13] ;
assign \14/3 = p_prod[5][12] ;
assign \14/4 = p_prod[6][11] ;
assign \14/5 = p_prod[7][10] ;
assign \14/6 = p_prod[8][9] ;
assign \14/7 = p_prod[9][8] ;
assign \14/8 = p_prod[10][7] ;
assign \14/9 = p_prod[11][6] ;
assign \14/10 = p_prod[12][5] ;
assign \14/11 = p_prod[13][4] ;
assign \14/12 = p_prod[14][3] ;
assign \14/13 = p_prod[15][2] ;
assign \15/0 = p_prod[1][15] ;
assign \15/1 = p_prod[2][14] ;
assign \15/2 = p_prod[3][13] ;
assign \15/3 = p_prod[4][12] ;
assign \15/4 = p_prod[5][11] ;
assign \15/5 = p_prod[6][10] ;
assign \15/6 = p_prod[7][9] ;
assign \15/7 = p_prod[8][8] ;
assign \15/8 = p_prod[9][7] ;
assign \15/9 = p_prod[10][6] ;
assign \15/10 = p_prod[11][5] ;
assign \15/11 = p_prod[12][4] ;
assign \15/12 = p_prod[13][3] ;
assign \15/13 = p_prod[14][2] ;
assign \15/14 = p_prod[15][1] ;
assign \16/0 = p_prod[0][15] ;
assign \16/1 = p_prod[1][14] ;
assign \16/2 = p_prod[2][13] ;
assign \16/3 = p_prod[3][12] ;
assign \16/4 = p_prod[4][11] ;
assign \16/5 = p_prod[5][10] ;
assign \16/6 = p_prod[6][9] ;
assign \16/7 = p_prod[7][8] ;
assign \16/8 = p_prod[8][7] ;
assign \16/9 = p_prod[9][6] ;
assign \16/10 = p_prod[10][5] ;
assign \16/11 = p_prod[11][4] ;
assign \16/12 = p_prod[12][3] ;
assign \16/13 = p_prod[13][2] ;
assign \16/14 = p_prod[14][1] ;
assign \16/15 = p_prod[15][0] ;
assign \17/0 = p_prod[0][14] ;
assign \17/1 = p_prod[1][13] ;
assign \17/2 = p_prod[2][12] ;
assign \17/3 = p_prod[3][11] ;
assign \17/4 = p_prod[4][10] ;
assign \17/5 = p_prod[5][9] ;
assign \17/6 = p_prod[6][8] ;
assign \17/7 = p_prod[7][7] ;
assign \17/8 = p_prod[8][6] ;
assign \17/9 = p_prod[9][5] ;
assign \17/10 = p_prod[10][4] ;
assign \17/11 = p_prod[11][3] ;
assign \17/12 = p_prod[12][2] ;
assign \17/13 = p_prod[13][1] ;
assign \17/14 = p_prod[14][0] ;
assign \18/0 = p_prod[0][13] ;
assign \18/1 = p_prod[1][12] ;
assign \18/2 = p_prod[2][11] ;
assign \18/3 = p_prod[3][10] ;
assign \18/4 = p_prod[4][9] ;
assign \18/5 = p_prod[5][8] ;
assign \18/6 = p_prod[6][7] ;
assign \18/7 = p_prod[7][6] ;
assign \18/8 = p_prod[8][5] ;
assign \18/9 = p_prod[9][4] ;
assign \18/10 = p_prod[10][3] ;
assign \18/11 = p_prod[11][2] ;
assign \18/12 = p_prod[12][1] ;
assign \18/13 = p_prod[13][0] ;
assign \19/0 = p_prod[0][12] ;
assign \19/1 = p_prod[1][11] ;
assign \19/2 = p_prod[2][10] ;
assign \19/3 = p_prod[3][9] ;
assign \19/4 = p_prod[4][8] ;
assign \19/5 = p_prod[5][7] ;
assign \19/6 = p_prod[6][6] ;
assign \19/7 = p_prod[7][5] ;
assign \19/8 = p_prod[8][4] ;
assign \19/9 = p_prod[9][3] ;
assign \19/10 = p_prod[10][2] ;
assign \19/11 = p_prod[11][1] ;
assign \19/12 = p_prod[12][0] ;
assign \20/0 = p_prod[0][11] ;
assign \20/1 = p_prod[1][10] ;
assign \20/2 = p_prod[2][9] ;
assign \20/3 = p_prod[3][8] ;
assign \20/4 = p_prod[4][7] ;
assign \20/5 = p_prod[5][6] ;
assign \20/6 = p_prod[6][5] ;
assign \20/7 = p_prod[7][4] ;
assign \20/8 = p_prod[8][3] ;
assign \20/9 = p_prod[9][2] ;
assign \20/10 = p_prod[10][1] ;
assign \20/11 = p_prod[11][0] ;
assign \21/0 = p_prod[0][10] ;
assign \21/1 = p_prod[1][9] ;
assign \21/2 = p_prod[2][8] ;
assign \21/3 = p_prod[3][7] ;
assign \21/4 = p_prod[4][6] ;
assign \21/5 = p_prod[5][5] ;
assign \21/6 = p_prod[6][4] ;
assign \21/7 = p_prod[7][3] ;
assign \21/8 = p_prod[8][2] ;
assign \21/9 = p_prod[9][1] ;
assign \21/10 = p_prod[10][0] ;
assign \22/0 = p_prod[0][9] ;
assign \22/1 = p_prod[1][8] ;
assign \22/2 = p_prod[2][7] ;
assign \22/3 = p_prod[3][6] ;
assign \22/4 = p_prod[4][5] ;
assign \22/5 = p_prod[5][4] ;
assign \22/6 = p_prod[6][3] ;
assign \22/7 = p_prod[7][2] ;
assign \22/8 = p_prod[8][1] ;
assign \22/9 = p_prod[9][0] ;
assign \23/0 = p_prod[0][8] ;
assign \23/1 = p_prod[1][7] ;
assign \23/2 = p_prod[2][6] ;
assign \23/3 = p_prod[3][5] ;
assign \23/4 = p_prod[4][4] ;
assign \23/5 = p_prod[5][3] ;
assign \23/6 = p_prod[6][2] ;
assign \23/7 = p_prod[7][1] ;
assign \23/8 = p_prod[8][0] ;
assign \24/0 = p_prod[0][7] ;
assign \24/1 = p_prod[1][6] ;
assign \24/2 = p_prod[2][5] ;
assign \24/3 = p_prod[3][4] ;
assign \24/4 = p_prod[4][3] ;
assign \24/5 = p_prod[5][2] ;
assign \24/6 = p_prod[6][1] ;
assign \24/7 = p_prod[7][0] ;
assign \25/0 = p_prod[0][6] ;
assign \25/1 = p_prod[1][5] ;
assign \25/2 = p_prod[2][4] ;
assign \25/3 = p_prod[3][3] ;
assign \25/4 = p_prod[4][2] ;
assign \25/5 = p_prod[5][1] ;
assign \25/6 = p_prod[6][0] ;
assign \26/0 = p_prod[0][5] ;
assign \26/1 = p_prod[1][4] ;
assign \26/2 = p_prod[2][3] ;
assign \26/3 = p_prod[3][2] ;
assign \26/4 = p_prod[4][1] ;
assign \26/5 = p_prod[5][0] ;
assign \27/0 = p_prod[0][4] ;
assign \27/1 = p_prod[1][3] ;
assign \27/2 = p_prod[2][2] ;
assign \27/3 = p_prod[3][1] ;
assign \27/4 = p_prod[4][0] ;
assign \28/0 = p_prod[0][3] ;
assign \28/1 = p_prod[1][2] ;
assign \28/2 = p_prod[2][1] ;
assign \28/3 = p_prod[3][0] ;
assign \29/0 = p_prod[0][2] ;
assign \29/1 = p_prod[1][1] ;
assign \29/2 = p_prod[2][0] ;
assign \30/0 = p_prod[0][1] ;
assign \30/1 = p_prod[1][0] ;
assign \31/0 = p_prod[0][0] ;
assign in1 = {1'b0,\1/0 ,\s76 ,\s126 ,\s158 ,\s159 ,\s180 ,\s181 ,\s182 ,\s183 ,\s195 ,\s196 ,\s197 ,\s198 ,\s199 ,\s200 ,\sf2 ,\sf3 ,\sf4 ,\sf5 ,\sf6 ,\sf7 ,\sf8 ,\sf9 ,\s201 ,\s194 ,\s179 ,\s157 ,\s125 ,\s75 ,\sf10 ,\31/0 };
assign in2 = {1'b0,\c76 ,\c126 ,\c158 ,\c159 ,\c180 ,\c181 ,\c182 ,\c183 ,\c195 ,\c196 ,\c197 ,\c198 ,\c199 ,\c200 ,\cf2 ,\cf3 ,\cf4 ,\cf5 ,\cf6 ,\cf7 ,\cf8 ,\cf9 ,\c201 ,1'b0,1'b0,1'b0,1'b0,1'b0,\cf10 ,1'b0,1'b0};

fullad csa0(\3/0 , \3/1 , \3/2 , \s1 , \c1 );
fullad csa1(\4/0 , \4/1 , \4/2 , \s2 , \c2 );
fullad csa2(\5/0 , \5/1 , \5/2 , \s3 , \c3 );
fullad csa3(\6/0 , \6/1 , \6/2 , \s4 , \c4 );
fullad csa4(\6/3 , \6/4 , \6/5 , \s5 , \c5 );
fullad csa5(\7/0 , \7/1 , \7/2 , \s6 , \c6 );
fullad csa6(\7/3 , \7/4 , \7/5 , \s7 , \c7 );
fullad csa7(\8/0 , \8/1 , \8/2 , \s8 , \c8 );
fullad csa8(\8/3 , \8/4 , \8/5 , \s9 , \c9 );
fullad csa9(\9/0 , \9/1 , \9/2 , \s10 , \c10 );
fullad csa10(\9/3 , \9/4 , \9/5 , \s11 , \c11 );
fullad csa11(\9/6 , \9/7 , \9/8 , \s12 , \c12 );
fullad csa12(\10/0 , \10/1 , \10/2 , \s13 , \c13 );
fullad csa13(\10/3 , \10/4 , \10/5 , \s14 , \c14 );
fullad csa14(\10/6 , \10/7 , \10/8 , \s15 , \c15 );
fullad csa15(\11/0 , \11/1 , \11/2 , \s16 , \c16 );
fullad csa16(\11/3 , \11/4 , \11/5 , \s17 , \c17 );
fullad csa17(\11/6 , \11/7 , \11/8 , \s18 , \c18 );
fullad csa18(\12/0 , \12/1 , \12/2 , \s19 , \c19 );
fullad csa19(\12/3 , \12/4 , \12/5 , \s20 , \c20 );
fullad csa20(\12/6 , \12/7 , \12/8 , \s21 , \c21 );
fullad csa21(\12/9 , \12/10 , \12/11 , \s22 , \c22 );
fullad csa22(\13/0 , \13/1 , \13/2 , \s23 , \c23 );
fullad csa23(\13/3 , \13/4 , \13/5 , \s24 , \c24 );
fullad csa24(\13/6 , \13/7 , \13/8 , \s25 , \c25 );
fullad csa25(\13/9 , \13/10 , \13/11 , \s26 , \c26 );
fullad csa26(\14/0 , \14/1 , \14/2 , \s27 , \c27 );
fullad csa27(\14/3 , \14/4 , \14/5 , \s28 , \c28 );
fullad csa28(\14/6 , \14/7 , \14/8 , \s29 , \c29 );
fullad csa29(\14/9 , \14/10 , \14/11 , \s30 , \c30 );
fullad csa30(\15/0 , \15/1 , \15/2 , \s31 , \c31 );
fullad csa31(\15/3 , \15/4 , \15/5 , \s32 , \c32 );
fullad csa32(\15/6 , \15/7 , \15/8 , \s33 , \c33 );
fullad csa33(\15/9 , \15/10 , \15/11 , \s34 , \c34 );
fullad csa34(\15/12 , \15/13 , \15/14 , \s35 , \c35 );
fullad csa35(\16/0 , \16/1 , \16/2 , \s36 , \c36 );
fullad csa36(\16/3 , \16/4 , \16/5 , \s37 , \c37 );
fullad csa37(\16/6 , \16/7 , \16/8 , \s38 , \c38 );
fullad csa38(\16/9 , \16/10 , \16/11 , \s39 , \c39 );
fullad csa39(\16/12 , \16/13 , \16/14 , \s40 , \c40 );
fullad csa40(\17/0 , \17/1 , \17/2 , \s41 , \c41 );
fullad csa41(\17/3 , \17/4 , \17/5 , \s42 , \c42 );
fullad csa42(\17/6 , \17/7 , \17/8 , \s43 , \c43 );
fullad csa43(\17/9 , \17/10 , \17/11 , \s44 , \c44 );
fullad csa44(\17/12 , \17/13 , \17/14 , \s45 , \c45 );
fullad csa45(\18/0 , \18/1 , \18/2 , \s46 , \c46 );
fullad csa46(\18/3 , \18/4 , \18/5 , \s47 , \c47 );
fullad csa47(\18/6 , \18/7 , \18/8 , \s48 , \c48 );
fullad csa48(\18/9 , \18/10 , \18/11 , \s49 , \c49 );
fullad csa49(\19/0 , \19/1 , \19/2 , \s50 , \c50 );
fullad csa50(\19/3 , \19/4 , \19/5 , \s51 , \c51 );
fullad csa51(\19/6 , \19/7 , \19/8 , \s52 , \c52 );
fullad csa52(\19/9 , \19/10 , \19/11 , \s53 , \c53 );
fullad csa53(\20/0 , \20/1 , \20/2 , \s54 , \c54 );
fullad csa54(\20/3 , \20/4 , \20/5 , \s55 , \c55 );
fullad csa55(\20/6 , \20/7 , \20/8 , \s56 , \c56 );
fullad csa56(\20/9 , \20/10 , \20/11 , \s57 , \c57 );
fullad csa57(\21/0 , \21/1 , \21/2 , \s58 , \c58 );
fullad csa58(\21/3 , \21/4 , \21/5 , \s59 , \c59 );
fullad csa59(\21/6 , \21/7 , \21/8 , \s60 , \c60 );
fullad csa60(\22/0 , \22/1 , \22/2 , \s61 , \c61 );
fullad csa61(\22/3 , \22/4 , \22/5 , \s62 , \c62 );
fullad csa62(\22/6 , \22/7 , \22/8 , \s63 , \c63 );
fullad csa63(\23/0 , \23/1 , \23/2 , \s64 , \c64 );
fullad csa64(\23/3 , \23/4 , \23/5 , \s65 , \c65 );
fullad csa65(\23/6 , \23/7 , \23/8 , \s66 , \c66 );
fullad csa66(\24/0 , \24/1 , \24/2 , \s67 , \c67 );
fullad csa67(\24/3 , \24/4 , \24/5 , \s68 , \c68 );
fullad csa68(\25/0 , \25/1 , \25/2 , \s69 , \c69 );
fullad csa69(\25/3 , \25/4 , \25/5 , \s70 , \c70 );
fullad csa70(\26/0 , \26/1 , \26/2 , \s71 , \c71 );
fullad csa71(\26/3 , \26/4 , \26/5 , \s72 , \c72 );
fullad csa72(\27/0 , \27/1 , \27/2 , \s73 , \c73 );
fullad csa73(\28/0 , \28/1 , \28/2 , \s74 , \c74 );
fullad csa74(\29/0 , \29/1 , \29/2 , \s75 , \c75 );
fullad csa75(\2/0 , \2/1 , \c1 , \s76 , \c76 );
fullad csa76(\4/3 , \s2 , \c3 , \s77 , \c77 );
fullad csa77(\5/3 , \5/4 , \s3 , \s78 , \c78 );
fullad csa78(\s4 , \s5 , \c6 , \s79 , \c79 );
fullad csa79(\7/6 , \s6 , \s7 , \s80 , \c80 );
fullad csa80(\8/6 , \8/7 , \s8 , \s81 , \c81 );
fullad csa81(\s9 , \c10 , \c11 , \s82 , \c82 );
fullad csa82(\s10 , \s11 , \s12 , \s83 , \c83 );
fullad csa83(\c13 , \c14 , \c15 , \s84 , \c84 );
fullad csa84(\10/9 , \s13 , \s14 , \s85 , \c85 );
fullad csa85(\s15 , \c16 , \c17 , \s86 , \c86 );
fullad csa86(\11/9 , \11/10 , \s16 , \s87 , \c87 );
fullad csa87(\s17 , \s18 , \c19 , \s88 , \c88 );
fullad csa88(\c20 , \c21 , \c22 , \s89 , \c89 );
fullad csa89(\s19 , \s20 , \s21 , \s90 , \c90 );
fullad csa90(\s22 , \c23 , \c24 , \s91 , \c91 );
fullad csa91(\13/12 , \s23 , \s24 , \s92 , \c92 );
fullad csa92(\s25 , \s26 , \c27 , \s93 , \c93 );
fullad csa93(\c28 , \c29 , \c30 , \s94 , \c94 );
fullad csa94(\14/12 , \14/13 , \s27 , \s95 , \c95 );
fullad csa95(\s28 , \s29 , \s30 , \s96 , \c96 );
fullad csa96(\c31 , \c32 , \c33 , \s97 , \c97 );
fullad csa97(\s31 , \s32 , \s33 , \s98 , \c98 );
fullad csa98(\s34 , \s35 , \c36 , \s99 , \c99 );
fullad csa99(\c37 , \c38 , \c39 , \s100 , \c100 );
fullad csa100(\16/15 , \s36 , \s37 , \s101 , \c101 );
fullad csa101(\s38 , \s39 , \s40 , \s102 , \c102 );
fullad csa102(\c41 , \c42 , \c43 , \s103 , \c103 );
fullad csa103(\s41 , \s42 , \s43 , \s104 , \c104 );
fullad csa104(\s44 , \s45 , \c46 , \s105 , \c105 );
fullad csa105(\c47 , \c48 , \c49 , \s106 , \c106 );
fullad csa106(\18/12 , \18/13 , \s46 , \s107 , \c107 );
fullad csa107(\s47 , \s48 , \s49 , \s108 , \c108 );
fullad csa108(\c50 , \c51 , \c52 , \s109 , \c109 );
fullad csa109(\19/12 , \s50 , \s51 , \s110 , \c110 );
fullad csa110(\s52 , \s53 , \c54 , \s111 , \c111 );
fullad csa111(\c55 , \c56 , \c57 , \s112 , \c112 );
fullad csa112(\s54 , \s55 , \s56 , \s113 , \c113 );
fullad csa113(\s57 , \c58 , \c59 , \s114 , \c114 );
fullad csa114(\21/9 , \21/10 , \s58 , \s115 , \c115 );
fullad csa115(\s59 , \s60 , \c61 , \s116 , \c116 );
fullad csa116(\22/9 , \s61 , \s62 , \s117 , \c117 );
fullad csa117(\s63 , \c64 , \c65 , \s118 , \c118 );
fullad csa118(\s64 , \s65 , \s66 , \s119 , \c119 );
fullad csa119(\24/6 , \24/7 , \s67 , \s120 , \c120 );
fullad csa120(\s68 , \c69 , \c70 , \s121 , \c121 );
fullad csa121(\25/6 , \s69 , \s70 , \s122 , \c122 );
fullad csa122(\s71 , \s72 , \c73 , \s123 , \c123 );
fullad csa123(\27/3 , \27/4 , \s73 , \s124 , \c124 );
fullad csa124(\28/3 , \s74 , \c75 , \s125 , \c125 );
fullad csa125(\s1 , \c2 , \c77 , \s126 , \c126 );
fullad csa126(\c4 , \c5 , \s78 , \s127 , \c127 );
fullad csa127(\c7 , \s79 , \c80 , \s128 , \c128 );
fullad csa128(\c8 , \c9 , \s80 , \s129 , \c129 );
fullad csa129(\c12 , \s81 , \s82 , \s130 , \c130 );
fullad csa130(\s83 , \s84 , \c85 , \s131 , \c131 );
fullad csa131(\c18 , \s85 , \s86 , \s132 , \c132 );
fullad csa132(\c87 , \c88 , \c89 , \s133 , \c133 );
fullad csa133(\s87 , \s88 , \s89 , \s134 , \c134 );
fullad csa134(\c25 , \c26 , \s90 , \s135 , \c135 );
fullad csa135(\s91 , \c92 , \c93 , \s136 , \c136 );
fullad csa136(\s92 , \s93 , \s94 , \s137 , \c137 );
fullad csa137(\c95 , \c96 , \c97 , \s138 , \c138 );
fullad csa138(\c34 , \c35 , \s95 , \s139 , \c139 );
fullad csa139(\s96 , \s97 , \c98 , \s140 , \c140 );
fullad csa140(\c40 , \s98 , \s99 , \s141 , \c141 );
fullad csa141(\s100 , \c101 , \c102 , \s142 , \c142 );
fullad csa142(\c44 , \c45 , \s101 , \s143 , \c143 );
fullad csa143(\s102 , \s103 , \c104 , \s144 , \c144 );
fullad csa144(\s104 , \s105 , \s106 , \s145 , \c145 );
fullad csa145(\c107 , \c108 , \c109 , \s146 , \c146 );
fullad csa146(\c53 , \s107 , \s108 , \s147 , \c147 );
fullad csa147(\s109 , \c110 , \c111 , \s148 , \c148 );
fullad csa148(\s110 , \s111 , \s112 , \s149 , \c149 );
fullad csa149(\c60 , \s113 , \s114 , \s150 , \c150 );
fullad csa150(\c62 , \c63 , \s115 , \s151 , \c151 );
fullad csa151(\s116 , \c117 , \c118 , \s152 , \c152 );
fullad csa152(\c66 , \s117 , \s118 , \s153 , \c153 );
fullad csa153(\c67 , \c68 , \s119 , \s154 , \c154 );
fullad csa154(\s120 , \s121 , \c122 , \s155 , \c155 );
fullad csa155(\c71 , \c72 , \s122 , \s156 , \c156 );
fullad csa156(\c74 , \s124 , \c125 , \s157 , \c157 );
fullad csa157(\s77 , \c78 , \c127 , \s158 , \c158 );
fullad csa158(\c79 , \s127 , \c128 , \s159 , \c159 );
fullad csa159(\c81 , \c82 , \s129 , \s160 , \c160 );
fullad csa160(\c83 , \c84 , \s130 , \s161 , \c161 );
fullad csa161(\c86 , \s131 , \c132 , \s162 , \c162 );
fullad csa162(\s132 , \s133 , \c134 , \s163 , \c163 );
fullad csa163(\c90 , \c91 , \s134 , \s164 , \c164 );
fullad csa164(\c94 , \s135 , \s136 , \s165 , \c165 );
fullad csa165(\s137 , \s138 , \c139 , \s166 , \c166 );
fullad csa166(\c99 , \c100 , \s139 , \s167 , \c167 );
fullad csa167(\s140 , \c141 , \c142 , \s168 , \c168 );
fullad csa168(\c103 , \s141 , \s142 , \s169 , \c169 );
halfad ha0(\c144 , \s169 , \sf1 , \cf1 );
fullad csa169(\c105 , \c106 , \s143 , \s170 , \c170 );
fullad csa170(\s144 , \c145 , \c146 , \s171 , \c171 );
fullad csa171(\s145 , \s146 , \c147 , \s172 , \c172 );
fullad csa172(\c112 , \s147 , \s148 , \s173 , \c173 );
fullad csa173(\c113 , \c114 , \s149 , \s174 , \c174 );
fullad csa174(\c115 , \c116 , \s150 , \s175 , \c175 );
fullad csa175(\s151 , \s152 , \c153 , \s176 , \c176 );
fullad csa176(\c119 , \s153 , \c154 , \s177 , \c177 );
fullad csa177(\c120 , \c121 , \s154 , \s178 , \c178 );
fullad csa178(\s123 , \c124 , \c157 , \s179 , \c179 );
fullad csa179(\s128 , \c129 , \c160 , \s180 , \c180 );
fullad csa180(\c130 , \s160 , \c161 , \s181 , \c181 );
fullad csa181(\c131 , \s161 , \c162 , \s182 , \c182 );
fullad csa182(\c133 , \s162 , \c163 , \s183 , \c183 );
fullad csa183(\c135 , \c136 , \s164 , \s184 , \c184 );
fullad csa184(\c137 , \c138 , \s165 , \s185 , \c185 );
fullad csa185(\c140 , \s166 , \c167 , \s186 , \c186 );
fullad csa186(\s167 , \s168 , \c169 , \s187 , \c187 );
fullad csa187(\c143 , \sf1 , \c170 , \s188 , \c188 );
fullad csa188(\s170 , \s171 , \c172 , \s189 , \c189 );
fullad csa189(\c148 , \s172 , \c173 , \s190 , \c190 );
fullad csa190(\c149 , \s173 , \c174 , \s191 , \c191 );
fullad csa191(\c150 , \s174 , \c175 , \s192 , \c192 );
fullad csa192(\c151 , \c152 , \s175 , \s193 , \c193 );
fullad csa193(\c123 , \s156 , \c179 , \s194 , \c194 );
fullad csa194(\s163 , \c164 , \c184 , \s195 , \c195 );
fullad csa195(\c165 , \s184 , \c185 , \s196 , \c196 );
fullad csa196(\c166 , \s185 , \c186 , \s197 , \c197 );
fullad csa197(\c168 , \s186 , \c187 , \s198 , \c198 );
fullad csa198(\cf1 , \s187 , \c188 , \s199 , \c199 );
fullad csa199(\c171 , \s188 , \c189 , \s200 , \c200 );
halfad ha1(\s189 , \c190 , \sf2 , \cf2 );
halfad ha2(\s190 , \c191 , \sf3 , \cf3 );
halfad ha3(\s191 , \c192 , \sf4 , \cf4 );
halfad ha4(\s192 , \c193 , \sf5 , \cf5 );
halfad ha5(\c176 , \s193 , \sf6 , \cf6 );
halfad ha6(\s176 , \c177 , \sf7 , \cf7 );
halfad ha7(\s177 , \c178 , \sf8 , \cf8 );
halfad ha8(\c155 , \s178 , \sf9 , \cf9 );
fullad csa200(\s155 , \c156 , \c194 , \s201 , \c201 );
halfad ha9(\30/0 , \30/1 , \sf10 , \cf10 );
halfad ha10(\s75 , \cf10 , \sf11 , \cf11 );
halfad ha11(\s125 , \cf11 , \sf12 , \cf12 );
halfad ha12(\s157 , \cf12 , \sf13 , \cf13 );
halfad ha13(\s179 , \cf13 , \sf14 , \cf14 );
halfad ha14(\s194 , \cf14 , \sf15 , \cf15 );
halfad ha15(\s201 , \cf15 , \sf16 , \cf16 );
fullad csa201(\sf9 , \c201 , \cf16 , \s202 , \c202 );
fullad csa202(\sf8 , \cf9 , \c202 , \s203 , \c203 );
fullad csa203(\sf7 , \cf8 , \c203 , \s204 , \c204 );
fullad csa204(\sf6 , \cf7 , \c204 , \s205 , \c205 );
fullad csa205(\sf5 , \cf6 , \c205 , \s206 , \c206 );
fullad csa206(\sf4 , \cf5 , \c206 , \s207 , \c207 );
fullad csa207(\sf3 , \cf4 , \c207 , \s208 , \c208 );
fullad csa208(\sf2 , \cf3 , \c208 , \s209 , \c209 );
fullad csa209(\s200 , \cf2 , \c209 , \s210 , \c210 );
fullad csa210(\s199 , \c200 , \c210 , \s211 , \c211 );
fullad csa211(\s198 , \c199 , \c211 , \s212 , \c212 );
fullad csa212(\s197 , \c198 , \c212 , \s213 , \c213 );
fullad csa213(\s196 , \c197 , \c213 , \s214 , \c214 );
fullad csa214(\s195 , \c196 , \c214 , \s215 , \c215 );
fullad csa215(\s183 , \c195 , \c215 , \s216 , \c216 );
fullad csa216(\s182 , \c183 , \c216 , \s217 , \c217 );
fullad csa217(\s181 , \c182 , \c217 , \s218 , \c218 );
fullad csa218(\s180 , \c181 , \c218 , \s219 , \c219 );
fullad csa219(\s159 , \c180 , \c219 , \s220 , \c220 );
fullad csa220(\s158 , \c159 , \c220 , \s221 , \c221 );
fullad csa221(\s126 , \c158 , \c221 , \s222 , \c222 );
fullad csa222(\s76 , \c126 , \c222 , \s223 , \c223 );
fullad csa223(\1/0 , \c76 , \c223 , \s224 , \c224 );


csa32 finaladd(in1, in2, out, ov);


endmodule